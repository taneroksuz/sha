import sha_const::*;

module sha_array(
  output logic [31 : 0] K_256 [0:63],
  output logic [63 : 0] K_512 [0:79],
  output logic [31 : 0] H_1 [0:4],
  output logic [31 : 0] H_224 [0:7],
  output logic [31 : 0] H_256 [0:7],
  output logic [63 : 0] H_384 [0:7],
  output logic [63 : 0] H_512 [0:7],
  output logic [63 : 0] H_512_224 [0:7],
  output logic [63 : 0] H_512_256 [0:7]
);
  timeunit 1ns;
  timeprecision 1ps;

  logic [31 : 0] k_256 [0:63];
  logic [63 : 0] k_512 [0:79];
  logic [31 : 0] h_1 [0:4];
  logic [31 : 0] h_224 [0:7];
  logic [31 : 0] h_256 [0:7];
  logic [63 : 0] h_384 [0:7];
  logic [63 : 0] h_512 [0:7];
  logic [63 : 0] h_512_224 [0:7];
  logic [63 : 0] h_512_256 [0:7];

  initial begin
    k_256[0]=32'h428a2f98; k_256[1]=32'h71374491; k_256[2]=32'hb5c0fbcf; k_256[3]=32'he9b5dba5; k_256[4]=32'h3956c25b; k_256[5]=32'h59f111f1; k_256[6]=32'h923f82a4; k_256[7]=32'hab1c5ed5;
    k_256[8]=32'hd807aa98; k_256[9]=32'h12835b01; k_256[10]=32'h243185be; k_256[11]=32'h550c7dc3; k_256[12]=32'h72be5d74; k_256[13]=32'h80deb1fe; k_256[14]=32'h9bdc06a7; k_256[15]=32'hc19bf174;
    k_256[16]=32'he49b69c1; k_256[17]=32'hefbe4786; k_256[18]=32'h0fc19dc6; k_256[19]=32'h240ca1cc; k_256[20]=32'h2de92c6f; k_256[21]=32'h4a7484aa; k_256[22]=32'h5cb0a9dc; k_256[23]=32'h76f988da;
    k_256[24]=32'h983e5152; k_256[25]=32'ha831c66d; k_256[26]=32'hb00327c8; k_256[27]=32'hbf597fc7; k_256[28]=32'hc6e00bf3; k_256[29]=32'hd5a79147; k_256[30]=32'h06ca6351; k_256[31]=32'h14292967;
    k_256[32]=32'h27b70a85; k_256[33]=32'h2e1b2138; k_256[34]=32'h4d2c6dfc; k_256[35]=32'h53380d13; k_256[36]=32'h650a7354; k_256[37]=32'h766a0abb; k_256[38]=32'h81c2c92e; k_256[39]=32'h92722c85;
    k_256[40]=32'ha2bfe8a1; k_256[41]=32'ha81a664b; k_256[42]=32'hc24b8b70; k_256[43]=32'hc76c51a3; k_256[44]=32'hd192e819; k_256[45]=32'hd6990624; k_256[46]=32'hf40e3585; k_256[47]=32'h106aa070;
    k_256[48]=32'h19a4c116; k_256[49]=32'h1e376c08; k_256[50]=32'h2748774c; k_256[51]=32'h34b0bcb5; k_256[52]=32'h391c0cb3; k_256[53]=32'h4ed8aa4a; k_256[54]=32'h5b9cca4f; k_256[55]=32'h682e6ff3;
    k_256[56]=32'h748f82ee; k_256[57]=32'h78a5636f; k_256[58]=32'h84c87814; k_256[59]=32'h8cc70208; k_256[60]=32'h90befffa; k_256[61]=32'ha4506ceb; k_256[62]=32'hbef9a3f7; k_256[63]=32'hc67178f2;

    k_512[0]=64'h428a2f98d728ae22; k_512[1]=64'h7137449123ef65cd; k_512[2]=64'hb5c0fbcfec4d3b2f; k_512[3]=64'he9b5dba58189dbbc; k_512[4]=64'h3956c25bf348b538;
    k_512[5]=64'h59f111f1b605d019; k_512[6]=64'h923f82a4af194f9b; k_512[7]=64'hab1c5ed5da6d8118; k_512[8]=64'hd807aa98a3030242; k_512[9]=64'h12835b0145706fbe;
    k_512[10]=64'h243185be4ee4b28c; k_512[11]=64'h550c7dc3d5ffb4e2; k_512[12]=64'h72be5d74f27b896f; k_512[13]=64'h80deb1fe3b1696b1; k_512[14]=64'h9bdc06a725c71235;
    k_512[15]=64'hc19bf174cf692694; k_512[16]=64'he49b69c19ef14ad2; k_512[17]=64'hefbe4786384f25e3; k_512[18]=64'h0fc19dc68b8cd5b5; k_512[19]=64'h240ca1cc77ac9c65;
    k_512[20]=64'h2de92c6f592b0275; k_512[21]=64'h4a7484aa6ea6e483; k_512[22]=64'h5cb0a9dcbd41fbd4; k_512[23]=64'h76f988da831153b5; k_512[24]=64'h983e5152ee66dfab;
    k_512[25]=64'ha831c66d2db43210; k_512[26]=64'hb00327c898fb213f; k_512[27]=64'hbf597fc7beef0ee4; k_512[28]=64'hc6e00bf33da88fc2; k_512[29]=64'hd5a79147930aa725;
    k_512[30]=64'h06ca6351e003826f; k_512[31]=64'h142929670a0e6e70; k_512[32]=64'h27b70a8546d22ffc; k_512[33]=64'h2e1b21385c26c926; k_512[34]=64'h4d2c6dfc5ac42aed;
    k_512[35]=64'h53380d139d95b3df; k_512[36]=64'h650a73548baf63de; k_512[37]=64'h766a0abb3c77b2a8; k_512[38]=64'h81c2c92e47edaee6; k_512[39]=64'h92722c851482353b;
    k_512[40]=64'ha2bfe8a14cf10364; k_512[41]=64'ha81a664bbc423001; k_512[42]=64'hc24b8b70d0f89791; k_512[43]=64'hc76c51a30654be30; k_512[44]=64'hd192e819d6ef5218;
    k_512[45]=64'hd69906245565a910; k_512[46]=64'hf40e35855771202a; k_512[47]=64'h106aa07032bbd1b8; k_512[48]=64'h19a4c116b8d2d0c8; k_512[49]=64'h1e376c085141ab53;
    k_512[50]=64'h2748774cdf8eeb99; k_512[51]=64'h34b0bcb5e19b48a8; k_512[52]=64'h391c0cb3c5c95a63; k_512[53]=64'h4ed8aa4ae3418acb; k_512[54]=64'h5b9cca4f7763e373;
    k_512[55]=64'h682e6ff3d6b2b8a3; k_512[56]=64'h748f82ee5defb2fc; k_512[57]=64'h78a5636f43172f60; k_512[58]=64'h84c87814a1f0ab72; k_512[59]=64'h8cc702081a6439ec;
    k_512[60]=64'h90befffa23631e28; k_512[61]=64'ha4506cebde82bde9; k_512[62]=64'hbef9a3f7b2c67915; k_512[63]=64'hc67178f2e372532b; k_512[64]=64'hca273eceea26619c;
    k_512[65]=64'hd186b8c721c0c207; k_512[66]=64'heada7dd6cde0eb1e; k_512[67]=64'hf57d4f7fee6ed178; k_512[68]=64'h06f067aa72176fba; k_512[69]=64'h0a637dc5a2c898a6;
    k_512[70]=64'h113f9804bef90dae; k_512[71]=64'h1b710b35131c471b; k_512[72]=64'h28db77f523047d84; k_512[73]=64'h32caab7b40c72493; k_512[74]=64'h3c9ebe0a15c9bebc;
    k_512[75]=64'h431d67c49c100d4c; k_512[76]=64'h4cc5d4becb3e42b6; k_512[77]=64'h597f299cfc657e2a; k_512[78]=64'h5fcb6fab3ad6faec; k_512[79]=64'h6c44198c4a475817;

    H_1[0]=32'h67452301; H_1[1]=32'hefcdab89; H_1[2]=32'h98badcfe; H_1[3]=32'h10325476; H_1[4]=32'hc3d2e1f0;

    H_224[0]=32'hc1059ed8; H_224[1]=32'h367cd507; H_224[2]=32'h3070dd17; H_224[3]=32'hf70e5939; H_224[4]=32'hffc00b31; H_224[5]=32'h68581511; H_224[6]=32'h64f98fa7; H_224[7]=32'hbefa4fa4;

    H_256[0]=32'h6a09e667; H_256[1]=32'hbb67ae85; H_256[2]=32'h3c6ef372; H_256[3]=32'ha54ff53a; H_256[4]=32'h510e527f; H_256[5]=32'h9b05688c; H_256[6]=32'h1f83d9ab; H_256[7]=32'h5be0cd19;

    H_384[0]=64'hcbbb9d5dc1059ed8; H_384[1]=64'h629a292a367cd507; H_384[2]=64'h9159015a3070dd17; H_384[3]=64'h152fecd8f70e5939; H_384[4]=64'h67332667ffc00b31; H_384[5]=64'h8eb44a8768581511; H_384[6]=64'hdb0c2e0d64f98fa7; H_384[7]=64'h47b5481dbefa4fa4;

    H_512[0]=64'h6a09e667f3bcc908; H_512[1]=64'hbb67ae8584caa73b; H_512[2]=64'h3c6ef372fe94f82b; H_512[3]=64'ha54ff53a5f1d36f1; H_512[4]=64'h510e527fade682d1; H_512[5]=64'h9b05688c2b3e6c1f; H_512[6]=64'h1f83d9abfb41bd6b; H_512[7]=64'h5be0cd19137e2179;

    H_512_224[0]=64'h8C3D37C819544DA2; H_512_224[1]=64'h73E1996689DCD4D6; H_512_224[2]=64'h1DFAB7AE32FF9C82; H_512_224[3]=64'h679DD514582F9FCF; H_512_224[4]=64'h0F6D2B697BD44DA8; H_512_224[5]=64'h77E36F7304C48942; H_512_224[6]=64'h3F9D85A86A1D36C8; H_512_224[7]=64'h1112E6AD91D692A1;

    H_512_256[0]=64'h22312194FC2BF72C; H_512_256[1]=64'h9F555FA3C84C64C2; H_512_256[2]=64'h2393B86B6F53B151; H_512_256[3]=64'h963877195940EABD; H_512_256[4]=64'h96283EE2A88EFFE3; H_512_256[5]=64'hBE5E1E2553863992; H_512_256[6]=64'h2B0199FC2C85B8AA; H_512_256[7]=64'h0EB72DDC81C52CA2;

  end

  assign K_256 = k_256;
  assign K_512 = k_512;
  assign H_1 = h_1;
  assign H_224 = h_224;
  assign H_256 = h_256;
  assign H_384 = h_384;
  assign H_512 = h_512;
  assign H_512_224 = h_512_224;
  assign H_512_256 = h_512_256;

endmodule
