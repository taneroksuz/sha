import sha_const::*;

module sha_block
(
  input logic rst,
  input logic clk
);
  timeunit 1ns;
  timeprecision 1ps;

endmodule
